--! 
--! \brief Version control file.
--! 
--! \author Gabriel Mariano Marcelino <gabriel.mm8@gmail.com>
--! 
--! \version 0.0.2
--! 
--! \date 2020/11/21
--! 

package version is

    constant GRISC_VERSION  : string := "0.0.2";

    constant GRISC_AUTHOR   : string := "Gabriel Mariano Marcelino";
    constant GRISC_EMAIL    : string := "gabriel.mm8@gmail.com";

    constant GRISC_STATUS   : string := "Development";

end version;
